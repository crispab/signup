# --- Constraints
constraint.required=Obligatorisk
constraint.min=Minvärde: {0}
constraint.max=Maxvärde: {0}
constraint.minLength=Minlängd: {0}
constraint.maxLength=Maxlängd: {0}
constraint.email=Epost

# --- Formats
format.date=Datum (''{0}'')
format.numeric=Numeriskt
format.real=Decimaltal

# --- Errors
error.invalid=Ogiltigt värde
error.invalid.java.util.Date=Ogiltigt datum
error.required=Obligatoriskt fält ej ifyllt
error.number=Fältet får bara innehålla siffror
error.real=Decimaltal förväntas
error.real.precision=Decimaltal med max {0} siffror inklusive {1} decimal(er) förväntas
error.min=Måste vara större än eller lika med {0}
error.min.strict=Måste vara större än {0}
error.max=Måste vara mindre än eller lika med {0}
error.max.strict=Måste vara mindre än {0}
error.minLength=Minlängd är {0}
error.maxLength=Maxlängd är {0}
error.email=Giltig epostadress förväntas
error.pattern=Måste uppfylla villkoret {0}
error.date=Giltigt datum förväntas

error.expected.date=Datum förväntas
error.expected.date.isoformat=Datum i ISO-format förväntas
error.expected.jodadate.format=Datum i JodaDate-format förväntas
error.expected.jsarray=Lista av värden förväntas
error.expected.jsboolean=Sant/falskt förväntas
error.expected.jsnumber=Tal förväntas
error.expected.jsobject=Objekt förväntas
error.expected.jsstring=Text förväntas
error.expected.jsnumberorjsstring=Text eller siffror förväntas
error.expected.keypathnode=Nod förväntas
error.expected.uuid=UUID förväntas

error.path.empty=Tom sökväg
error.path.missing=Sökväg saknas
error.path.result.multiple=Sökvägen ger fler än ett resultat
