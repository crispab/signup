# SignUp messages


# ----------------------------------------------
# Default messages in Play translated to Swedish

# --- Constraints
user.updateimage.standard.heading=Standardbild
constraint.required=Obligatorisk
constraint.min=Minvärde: {0}
constraint.max=Maxvärde: {0}
constraint.minLength=Minlängd: {0}
constraint.maxLength=Maxlängd: {0}
constraint.email=Epost

# --- Formats
format.date=Datum (''{0}'')
format.numeric=Numeriskt
format.real=Decimaltal

# --- Errors
error.invalid=Ogiltigt värde
error.invalid.java.util.Date=Ogiltigt datum
error.required=Obligatoriskt fält ej ifyllt
error.number=Fältet får bara innehålla siffror
error.real=Decimaltal förväntas
error.real.precision=Decimaltal med max {0} siffror inklusive {1} decimal(er) förväntas
error.min=Måste vara större än eller lika med {0}
error.min.strict=Måste vara större än {0}
error.max=Måste vara mindre än eller lika med {0}
error.max.strict=Måste vara mindre än {0}
error.minLength=Minlängd är {0}
error.maxLength=Maxlängd är {0}
error.email=Giltig epostadress förväntas
error.pattern=Måste uppfylla villkoret {0}
error.date=Giltigt datum förväntas

error.expected.date=Datum förväntas
error.expected.date.isoformat=Datum i ISO-format förväntas
error.expected.jodadate.format=Datum i JodaDate-format förväntas
error.expected.jsarray=Lista av värden förväntas
error.expected.jsboolean=Sant/falskt förväntas
error.expected.jsnumber=Tal förväntas
error.expected.jsobject=Objekt förväntas
error.expected.jsstring=Text förväntas
error.expected.jsnumberorjsstring=Text eller siffror förväntas
error.expected.keypathnode=Nod förväntas
error.expected.uuid=UUID förväntas

error.path.empty=Tom sökväg
error.path.missing=Sökväg saknas
error.path.result.multiple=Sökvägen ger fler än ett resultat
navigation.home=Hem
errorpage.oops=Oj! Nu blev det visst fel.
errorpage.details=Tekniska detaljer
errorpage.startpage=Till startsidan
index.welcome=Välkommen till {0}
index.description.1={0} är en tjänst för grupper som vill ha ordning på sina sammankomster.
index.description.2=Du kan lägga upp nya sammankomster i gruppens kalender och medlemmarna kan själva gå in och markera ifall de kan komma eller inte.
index.description.3={0} skickar inbjudningar och påminnelser till alla medlemmar i gruppen för varje sammankomst.
navigation.users=Användare
login.login=Logga in
login.failed=Felaktig epostadress eller lösenord.
login.google=Logga in med Google
login.facebook=Logga in med Facebook
page.navbar.showhide=Visa/dölj navigation
navigation.mypage=Min sida
navigation.logout=Logga ut
login.email=Epost
login.password=Lösenord
login.with.password=Logga in med lösenord
login.with.social=Logga in med sociala media
errorpage.title=Fel
http.notfound=Sidan du försökte gå till finns inte
http.error=Sidan du försökte gå till kan inte visas
http.badrequest=Sidan du försökte gå till kan inte visas
status.on=Kommer
status.off=Kommer inte
status.maybe=Kanske
status.unregistered=Har inte svarat
application.logout=Du har loggats ut!
error.application.authfail=Nädu, det här får du inte göra utan att logga in som administratör!
login.nonexistentemail=Det finns ingen användare med epostadressen: {0}
login.unknownerror=Okänt fel
login.socialfail=Det gick inte att logga in via {0}: {1}
error.signup.eventcancelled=Sammankomsten är inställd. Det går inte att anmäla sig.
participation.people={0} i sällskapet
participation.updated=Anmälan uppdaterad för {0}: {1}
user.reminder=En påminnelse om sammankomsten kommer att skickas till {0}
event.cancelled.noreminders=Sammankomsten är inställd. Det går inte att skicka påminnelser.
user.upload.nofile=Du måste välja en bild från datorn
user.upload.error=Något gick snett vid inläsningen. Prova en annan bild.
error.signup.email.alreadyinuse=Epostadressen används av någon annan
error.signup.password.toshort=Lösenordet måste vara minst 8 tecken!!!
mail.sentreminders={0} har skickat påminnelse till {1} medlem(mar)
mail.failedreminder=Misslyckades att skicka påminnelse till {0}. {1}: {2}
mail.sentonereminder={0} har skickat påminnelse till {1}
slack.failedreminder=Misslyckades att skicka chattmeddelande på Slack. {0}: {1}
slack.sentreminders={0} har skickat chattmeddelande på Slack
excel.signups=Anmälningar
excel.firsname=Förnamn
excel.lastname=Efternamn
excel.email=Epost
excel.status=Status
excel.people=Antal
excel.date=Datum
excel.guest.heading=Gäst?
excel.guest=Gäst
excel.late.heading=Sen?
excel.late=Sen
excel.comment=Kommentar
event.remindersent=En påminnelse om sammankomsten kommer att skickas till alla delatagare som inte redan meddelat sig.
event.createdby=Sammankomsten skapad av {0}
event.remindersent.all=En inbjudan till sammankomsten håller på att skickas till alla
event.cancelled.noedit=Sammankomsten är inställd. Det går inte att redigera. Skapa en ny istället.
event.cancelledby=Sammankomsten inställd av {0}. Orsak: {1}
error.signup.endtime=Sluttid måste vara efter starttid
error.signup.lastsignup=Sista anmälningsdag måste vara före själva sammankomsten
navigation.groups=Grupper
event.eventpassed=Denna sammankomst har redan inträffat!
event.signupdatepassed=Sista anmälningsdatum har passerats.
event.full=Sammankomsten är fullbokad. Prova att kontrollera vid ett senare tillfälle ifall någon plats blivit ledig.
event.time=Tid:
event.venue=Plats:
event.maxparticipants=Max antal deltagare:
event.fullybooked=(fullbokat)
event.lastsignup=Sista anmälningsdag {0}
calendar.google=Google
calendar.online=(online)
calendar.outlookcom=Outlook.com
calendar.yahoo=Yahoo
calendar.outlook=Outlook
calendar.apple=Apple Kalender
calendar.add=Lägg till i kalender
event.excel=Som Excel
event.reminders=Påminnelser
event.notifications=Händelser
event.guests=Gäster
event.noguests=Inga extra gäster
event.members=Medlemmar
event.actions=Åtgärder
event.edit=Redigera sammankomst
event.remind=Påminn de som inte svarat
event.cancel=Ställ in
edit.remove=Ta bort
event.numberof={0} st
event.reminder.heading=Vill du e-posta de som ännu inte svarat?
event.reminder.warning=Du håller på att skicka en påminnelse via e-post till alla inbjudna delatagare till sammankomsten {0} som ännu inte svarat.
edit.continue=Vill du fortsätta?
button.cancel=Avbryt
event.reminder.action=Skicka påminnelse
event.cancel.heading=Vill du ställa in sammankomsten?
event.cancel.warning=Du håller på att ställa in sammankomsten {0} och meddela alla deltagare.
event.cancel.reason=Orsak
button.abort=Avbryt
event.cancel.action=Ställ in
calendar.event=Sammankomst: {0}
event.edit.title=Redigera sammankomst {0}
edit.new=Ny
edit.edit=Redigera
event.new=Ny sammankomst
event.edit.name=Namn
event.edit.name.error=Fyll i ett namn på sammankomsten
event.edit.description.error=Beskrivning sakna
event.edit.description=Beskrivning
event.edit.venue=Plats
event.edit.venue.error=Fyll i en plats där sammankomsten äger rum
event.edit.date=Dag
event.edit.date.error=Ogiltigt datum eller klockslag
event.edit.time.from=från kl
event.edit.time.to=till kl
event.edit.last=Sista anmälningsdag
event.edit.sameday=samma dag, eller
event.edit.last.error=Sista anmälningsdag får inte vara efter sammankomsten
event.edit.invited=Hantering av inbjudna
event.edit.invitedonly=Bara inbjudna får komma
event.edit.allowextrafriends=Inbjudna får ta med extra vänner
edit.error=Inmatningsfel
event.edit.reminder=Påminnelse
event.edit.reminder.description=Två påminnelser kommer att göras helt automatiskt med början {0} dagar innan sammankomsten.
event.edit.reminder.checkbox=Skicka påminnelse/inbjudan till alla när jag sparar
event.edit.reminder.immediately=Det går även att begära att ett utskick görs direkt när sammankomsten skapas:
button.save=Spara
event.showcancelled.title=Sammankomsten är inställd.
event.remove.heading=Vill du ta bort sammankomsten?
event.remove.warning=Du håller på att ta bort sammankomsten {0}.
event.reminder.future=Påminnelse kommer automatiskt att skickas {0}
event.late.heading=Sen anmälan
event.late.text=Anmälde sig {0}, vilket är efter sista anmälningsdag.
event.removeguest.heading=Vill du ta bort gästen?
event.removeguest.warning=Du håller på att ta bort gästen {0} {1} från sammankomsten {2}.
event.addguest=Ny gäst
event.notify.cancelled=Inställd sammankomst:
event.cancel.reason.none=Ej angiven
event.notify.reminder=Dags att anmäla sig till sammankomsten
event.notify.updated=Uppdaterad anmälan i sammankomsten
participation.comment=Kommentar
event.notify.cancelledingroup=Inställt i gruppen {0}
event.notify.hello=Hej {0}!
event.notify.cancelled.message=Tyvärr har denna sammankomst blivit inställd.
event.notify.reminder.message=Nu är det dags att anmäla sig till nästa sammankomst.
event.notify.reminder.signup=Till anmälningssidan →
group.addgroup=Ny grupp
group.remove.heading=Vill du ta bort gruppen?
group.remove.warning=Du håller på att ta bort gruppen {0}.
navigation.events=Sammankomster
group.events.showfuture=Visa bara framtida
group.events.showall=Visa alla
group.event.cancelled=Inställt:
group.members=Medlemmar
group.members.count=({0} st)
group.member.remove.warning=Du håller på att ta bort medlemmen {0} {1}.
group.member.remove.heading=Vill du ta bort medlemmen?
group.addmember=Ny medlem
group.edit=Redigera grupp {0}
group.edit.name=Namn
group.edit.name.error=Fyll i ett namn på gruppen
group.edit.description=Beskrivning
group.edit.description.error=Det här var en underlig beskrivning
group.edit.email.title=Konfigurering av epost från gruppen
group.edit.email.sender=Avsändare
group.edit.email.sender.error=Fyll i adressen till den som skall stå som avsändare
group.edit.email.subjectprefix=Rubrikprefix
group.edit.email.subjectprefix.error=Fyll i vad mailrubriker skall börja med
navigation.membership=Ny medlem
group.new=Ny grupp
membership.heading=Ny medlem i {0}
membership.existinguser=Befintlig användare
option.noperson=Ingen vald
membership.error.selectuser=Välj en användare som medlem
membership.add=Lägg till
membership.new=Ny användare
participation.heading=Anmälan till {0}
navigation.participation=Anmälan
participation.remind=Påminn deltagaren
participation.reminder.heading=Vill du e-posta deltagaren?
participation.reminder.warning=Du håller på att skicka en påminnelse via e-post till {0} {1} om sammankomsten {2}.
participation.error.attendance=Välj om du kommer eller inte
participation.participants=Antal deltagare:
participation.save=Anmäl
participation.guest.heading=Ny gäst till {0}
navigation.guest=Ny gäst
participation.guest.error=Välj en användare som gäst
user.edit=Redigera användare {0} {1}
user.new=Ny användare
user.edit.firstname=Förnamn
user.edit.lastname=Efternamn
user.edit.firstname.error=Fyll i förnamn
user.edit.lastname.error=Fyll i efternamn
user.edit.email=Epost
user.edit.email.error=Fyll i en korrekt epostadress
user.edit.phone=Telefonnummer
user.edit.phone.error=Ogiltigt telefonnummer
user.edit.description=Beskrivning
user.edit.description.error=Va?? Skum beskrivning.
user.edit.password=Lösenord
user.edit.password.error=Du måste ange ett lösenord på minst 8 tecken
user.edit.adminperm=Har administratörsbehörighet
user.edit.role=Roll
user.role.administrator=Administratör
user.remove.heading=Vill du ta bort användaren?
user.remove.warning=Du håller på att ta bort användaren {0} {1}.
button.use=Använd
navigation.updateimage=Byt bild
user.updateimage.standard.row1=Om du har registrerat dig på 
user.updateimage.standard.row2=och kopplat en bild till din epostadress visas den bilden.
user.updateimage.standard.row3=Annars visas en anonym bild.
user.updateimage.own.heading=Egen bild
user.updateimage.own.row1=Välj en bild på datorn och använd den som profilbild.
user.updateimage.own.row2=Bilden kommer automatiskt att zoomas in på ansiktet, beskäras och skalas om.
user.updateimage=Byt bild för {0} {1} 
excel.description=Beskrivning
